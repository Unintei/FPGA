`timescale  1ns/1ns

////////////////////////////////////////////////////////////////////////

module  tb_PWM_Led();

//********************************************************************//
//****************** Parameter and Internal Signal *******************//
//********************************************************************//
//wire  define
wire    	[2:0]   	led_out     ;
wire		[5:0]		stear_s;
//reg   define
reg             sys_clk     ;
reg             sys_rst_n   ;

//********************************************************************//
//***************************** Main Code ****************************//
//********************************************************************//
//初始化系统时钟、全局复位
initial begin
	sys_clk    = 1'b1;
    sys_rst_n <= 1'b0;
    #20
	#1
    sys_rst_n <= 1'b1;
end

//sys_clk:模拟系统时钟，每10ns电平翻转一次，周期为20ns，频率为50Mhz
always #10 sys_clk = ~sys_clk;

//********************************************************************//
//*************************** Instantiation **************************//
//********************************************************************//
//-------------------- water_led_inst --------------------
PWM_Led   
#(
    .CNT_MAX    (26'd20000),
	.T_s		(15'd3)
	)
PWM_Led_inst
(
    .sys_clk    (sys_clk    ),  //input          sys_clk
    .sys_rst_n  (sys_rst_n  ),  //input          sys_rst_n
           
    .stear_s    (stear_s    ),   //output  [3:0]  led_out
	.led_out 	(led_out    )
); 	

endmodule
