/*****************************************************
	动态数码管 
	2023/11/21    1s切换一位
*****************************************************/
module  jsq
#(
//****************************************************//

//定义晶振频率50M
    parameter CNT_MAX = 26'd50_000_000 
	 
//****************************************************//
)
(
    input   wire            sys_clk     ,   //输入工作时钟,频率50MHz
    input   wire            sys_rst_n   ,   //输入复位信号,低电平有效

    output  wire            end_cnt0          //输出行同步信号

);

//reg   define
reg     [25:0]  cnt0         ;    //1s

//********************************************************************//
//***************************** Main Code ****************************//
//********************************************************************//

//cnt0:计数器计数1s
always @(posedge sys_clk or negedge sys_rst_n)begin
    if(!sys_rst_n)begin  
        cnt0 <= 0;
    end
    else if(add_cnt0)begin
        if(end_cnt0)
            cnt0 <= 0;   
        else
            cnt0 <= cnt0 + 1;
    end
end

assign add_cnt0 = 1;     //对时钟计数，计数条件始终有效
assign end_cnt0 = add_cnt0 && cnt0== CNT_MAX -1 ;//计数1s 

endmodule
