`timescale 1 ns/1 ns

module key_module_tb();

//parameter define
//Ϊ�����̷���ʱ�䣬���ǽ���������ʱ��ֵ��С
//��λ����Ȼ����Ͳ�������ֵ����һ��
//Ҳ���Խ���Щ����ֵ�ĳɺͲ�������ֵһ��
parameter   CNT_1MS  = 20'd19   ,
            CNT_11MS = 21'd69   ,
            CNT_41MS = 22'd149  ,
            CNT_51MS = 22'd199  ,
            CNT_60MS = 22'd249  ;

//wire  define
wire    [2:0]        key_vld    ;   //�����󰴼��ź�

//reg   define
reg             clk             ;   //����ʱ���ź�
reg             rst_n           ;   //���渴λ�ź�
reg     [2:0]    key_in         ;   //ģ�ⰴ������
reg     [21:0]  tb_cnt          ;   //ģ�ⰴ������������

//ʱ�����ڣ���λΪns�����ڴ��޸�ʱ�����ڡ�
parameter CYCLE    = 20;

//��λʱ�䣬��ʱ��ʾ��λ3��ʱ�����ڵ�ʱ�䡣
parameter RST_TIME = 3 ;

//�����Ե�ģ������
key_module  uut0(
    .clk         (clk      ), 
    .rst_n       (rst_n    ),
    .key_in      (key_in   ),
    .key_vld     (key_vld  )
);

initial begin
    clk    =1'b1;
    rst_n <=1'b0;
    key_in<=1'b0;
    #20
    rst_n <=1'b1;
end

//clkģ��ʱ�ӣ�50MHz
always #10 clk =~clk;

//tb_cnt:�������̼�������ͨ���ü������ļ���ʱ����ģ�ⰴ���Ķ�������
always@(posedge clk or negedge rst_n)
    if(rst_n == 1'b0)
        tb_cnt <= 22'b0;
    else    if(tb_cnt == CNT_60MS)
   //������������CNT_60MS���һ�ΰ����Ӱ��µ��ͷŵ���������
        tb_cnt <= 22'b0;
    else    
        tb_cnt <= tb_cnt + 1'b1;

//key_in:���������������ģ�ⰴ�����������
always@(posedge clk or negedge rst_n)
    if(rst_n == 1'b0)
        key_in <= 1'b1;     //����δ����ʱ��״̬ΪΪ�ߵ�ƽ
    else    if((tb_cnt >= CNT_1MS && tb_cnt <= CNT_11MS)
                || (tb_cnt >= CNT_41MS && tb_cnt <= CNT_51MS))
    //�ڸü��������ڲ����Ǹ������0��1��ģ��10ms��ǰ������10ms�ĺ󶶶�
        key_in <= {$random} % 2;    
    else    if(tb_cnt >= CNT_11MS && tb_cnt <= CNT_41MS)
        key_in <= 1'b0;
    //��������10ms��ǰ�������ȶ��ڵ͵�ƽ������ʱ�������CNT_MAX
    else
        key_in <= 1'b1;

endmodule

