module moduleRGB_Control(
	input	clk_RGB_Control,
	input	rst_n,
	input [7:0] uart_data,
	input	tx_done,		//一帧(24bit)数据结束标志，
	output	tx_en,			//发送数据使能
	output	reg	[23:0]	RGB
);

//-------------接口信号------------//
reg	[31:0]	cnt;
reg 	[4:0]	k;				
reg 	tx_en_r;                   // tx_en_r发送数据控制使能
reg   [23:0]	RGB_reg	[8:0] ;  //存RGB数据的数组
//--------------------------------//
//控制一帧（24bit）数据结束
//当复位时，清零
//否则，信号由RZ_Code模块输出tx_done提供
reg 	tx_done_r0;                
always @(posedge clk_RGB_Control or negedge rst_n) begin
	if(!rst_n)	begin
		tx_done_r0 <= 0;
	end
	else	begin
		tx_done_r0 <= tx_done;
	end
end

//--------------------------------//
//状态选择
reg [1:0]   mode_1 ;
reg [7:0]   mode_2 ;
reg         flag_1;
reg         flag_2;
reg [1:0]   time_flag_1 ;
reg [3:0]   time_flag_2 ;
reg [40:0]  Count1 ;
reg [40:0]  Count2 ; 
reg [32:0]  t ;
reg [9:0]   mode ;
//------------------------------------//


//----------------速度选择--------------------// t = 时间 * 5_000_0000
always @(posedge clk_RGB_Control)  begin
    if (uart_data[0])   begin  
        t <= 33'd4999_999 ; //  T = 0.1S  
	end
	else if (uart_data[1])   begin
        t <= 33'd4999_999*5 ;  //  T = 3S
	end
	else  begin
        t = 33'd49999_999 ;   // T =1S	 
	end
end

//-------------------------------//


//-----------模式控制模块-----------//
always @(posedge clk_RGB_Control)  begin
    if (uart_data[2])   begin
	    flag_1 <= 0 ;
	    flag_2 <= 1 ;							 
	end
	else if (uart_data[3])   begin    
	    flag_1 <= 1 ;
	    flag_2 <= 0 ;
	end
	else  begin     
        flag_1 <= 0 ;	
	    flag_2 <= 0 ;
	end	
end


//-------------时间控制模块计数器----------------------//
always @(posedge clk_RGB_Control) begin 
    if(flag_1) begin
        if(Count1 == t)      
           Count1 <= 0 ;
	    else 
           Count1 <= Count1 + 1 ; 
        end
    else
        Count1 <= 0 ;	
end

always @(posedge clk_RGB_Control) begin 
    if(flag_2) begin
		if(Count2 == 8 * (t+1))    
            Count2 <= 0 ;
		else 
            Count2 <= Count2 + 1 ;
		end	
	else                           
            Count2 <= 0 ;
end

//--------------状态模块----------------------//
always @(posedge clk_RGB_Control) begin
     if(Count1 == 0)                         time_flag_1 <= 2'd0 ;
	  else if(Count1 == 5)                   time_flag_1 <= 2'd1 ;
	  else if(Count1 == (t+1)/2)             time_flag_1 <= 2'd2 ;
  
end

always @(posedge clk_RGB_Control) begin
     if     (Count2 == 0)                   time_flag_2 <= 16'd0 ;
  
	  else if(Count2 == 10)                  time_flag_2 <= 16'd1 ;
	  
	  else if(Count2 == t)                   time_flag_2 <= 16'd2 ;
	  
	  else if(Count2 == 2 * (t+1)-1)         time_flag_2 <= 16'd3 ; 
	  
     else if(Count2 == 3 * (t+1)-1)         time_flag_2 <= 16'd4 ; 
	  
	  else if(Count2 == 4 * (t+1)-1)         time_flag_2 <= 16'd5 ; 
	   
	  else if(Count2 == 5 * (t+1)-1)         time_flag_2 <= 16'd6 ;
	  
	  else if(Count2 == 6 * (t+1)-1)         time_flag_2 <= 16'd7 ; 
	  
	  else if(Count2 == 7 * (t+1)-1)         time_flag_2 <= 16'd8 ; 
  
end

//----------模式的状态变化----------//
always @(*) begin
     if     (time_flag_1 == 2'd0)    mode_1 <= 2'b00 ;

	  else if(time_flag_1 == 2'd1)    mode_1 <= 2'b01 ;
	  
	  else if(time_flag_1 == 2'd2)    mode_1 <= 2'b10 ;
 
end



always @(posedge clk_RGB_Control) begin
     if     (time_flag_2 == 16'd0)   mode_2 <= 8'b00000000 ;
   
	  else if(time_flag_2 == 16'd1)   mode_2 <= 8'b00000001 ;
	  
	  else if(time_flag_2 == 16'd2)   mode_2 <= 8'b00000010 ; 
	  
	  else if(time_flag_2 == 16'd3)   mode_2 <= 8'b00000100 ; 
	  
     else if(time_flag_2 == 16'd4)   mode_2 <= 8'b00001000 ; 
	  
	  else if(time_flag_2 == 16'd5)   mode_2 <= 8'b00010000 ; 
	  
	  else if(time_flag_2 == 16'd6)   mode_2 <= 8'b00100000 ;  
	  
	  else if(time_flag_2 == 16'd7)   mode_2 <= 8'b01000000 ; 
	  
	  else if(time_flag_2 == 16'd8)   mode_2 <= 8'b10000000 ; 
  
end

always @(posedge clk_RGB_Control) begin
    mode <= {mode_2, mode_1} ;
	if(uart_data[4])begin
//1. 闪烁+绿色单色移位循环
// 如果count1等于多少多少的时候，RGB_reg等于多少多少，就达到了固定时间切换状态的效果
    case(mode)    
	   10'b0000000001 :  begin
	   RGB_reg	[0]	<= 24'b00000000_11111110_00000000; // 红
		RGB_reg	[1]	<= 24'b11001101_11111110_00000000; // 橙
		RGB_reg	[2]	<= 24'b11111110_11111110_00000000; // 黄
		RGB_reg	[3]	<= 24'b11111110_00000000_00000000; // 绿
		RGB_reg	[4]	<= 24'b11111110_00000000_11111110; // 青
		RGB_reg	[5]	<= 24'b00000000_00000000_11111110; // 蓝
		RGB_reg	[6]	<= 24'b00000000_11001100_11001100; // 紫
		RGB_reg	[7]	<= 24'b11111110_11111110_11111110; // 白
		RGB_reg	[8]	<= 24'b11111111_11111111_11111111;
		end

      10'b0000000010 :  begin
	  	RGB_reg	[0]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[1]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[2]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[3]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[4]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[5]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[6]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[7]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[8]	<= 24'b00000000_00000000_00000000;
		end
		
		// 绿色单色移位循环
		10'b0000000100 :  begin
	  	RGB_reg	[0]	<= 24'b11111110_00000000_00000000; 
		RGB_reg	[1]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[2]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[3]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[4]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[5]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[6]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[7]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[8]	<= 24'b00000000_00000000_00000000;
		end
		
		10'b0000001000 :  begin
	  	RGB_reg	[0]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[1]	<= 24'b11111110_00000000_00000000; 
		RGB_reg	[2]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[3]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[4]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[5]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[6]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[7]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[8]	<= 24'b00000000_00000000_00000000;
		end
		
		10'b0000010000 :  begin
	  	RGB_reg	[0]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[1]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[2]	<= 24'b11111110_00000000_00000000; 
		RGB_reg	[3]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[4]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[5]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[6]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[7]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[8]	<= 24'b00000000_00000000_00000000;
		end
		
		10'b0000100000 :  begin
	  	RGB_reg	[0]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[1]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[2]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[3]	<= 24'b11111110_00000000_00000000; 
		RGB_reg	[4]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[5]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[6]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[7]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[8]	<= 24'b00000000_00000000_00000000;
		end
		
		10'b0001000000 :  begin
	  	RGB_reg	[0]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[1]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[2]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[3]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[4]	<= 24'b11111110_00000000_00000000; 
		RGB_reg	[5]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[6]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[7]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[8]	<= 24'b00000000_00000000_00000000;
		end
		
		10'b0010000000 :  begin
	  	RGB_reg	[0]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[1]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[2]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[3]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[4]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[5]	<= 24'b11111110_00000000_00000000; 
		RGB_reg	[6]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[7]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[8]	<= 24'b00000000_00000000_00000000;
		end
		
		10'b0100000000 :  begin
	  	RGB_reg	[0]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[1]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[2]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[3]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[4]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[5]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[6]	<= 24'b11111110_00000000_00000000; 
		RGB_reg	[7]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[8]	<= 24'b00000000_00000000_00000000;
		end
		
		10'b1000000000 :  begin
	  	RGB_reg	[0]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[1]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[2]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[3]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[4]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[5]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[6]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[7]	<= 24'b11111110_00000000_00000000; 
		RGB_reg	[8]	<= 24'b00000000_00000000_00000000; // 白
		end
		endcase
	end
	else if(uart_data[5]) begin  
//2. 闪烁+七彩色移位循环 
	case(mode)    
	   10'b0000000001 :  begin
	   RGB_reg	[0]	<= 24'b00000000_11111110_00000000; // 红
		RGB_reg	[1]	<= 24'b11001101_11111110_00000000; // 橙
		RGB_reg	[2]	<= 24'b11111110_11111110_00000000; // 黄
		RGB_reg	[3]	<= 24'b11111110_00000000_00000000; // 绿
		RGB_reg	[4]	<= 24'b11111110_00000000_11111110; // 青
		RGB_reg	[5]	<= 24'b00000000_00000000_11111110; // 蓝
		RGB_reg	[6]	<= 24'b00000000_11001100_11001100; // 紫
		RGB_reg	[7]	<= 24'b11111110_11111110_11111110; // 白
		RGB_reg	[8]	<= 24'b11111111_11111111_11111111;
		end

      10'b0000000010 :  begin
	  	RGB_reg	[0]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[1]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[2]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[3]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[4]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[5]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[6]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[7]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[8]	<= 24'b00000000_00000000_00000000;
		end

      //红绿蓝白红绿蓝白循环
		10'b0000000100 :  begin
	   RGB_reg	[0]	<= 24'b00000000_11111110_00000000; // 红
		RGB_reg	[1]	<= 24'b11001101_11111110_00000000; // 橙
		RGB_reg	[2]	<= 24'b11111110_11111110_00000000; // 黄
		RGB_reg	[3]	<= 24'b11111110_00000000_00000000; // 绿
		RGB_reg	[4]	<= 24'b11111110_00000000_11111110; // 青
		RGB_reg	[5]	<= 24'b00000000_00000000_11111110; // 蓝
		RGB_reg	[6]	<= 24'b00000000_11001100_11001100; // 紫
		RGB_reg	[7]	<= 24'b11111110_11111110_11111110; // 白
		RGB_reg	[8]	<= 24'b11111111_11111111_11111111;
		end
		
		10'b0000001000 :  begin
	  	RGB_reg	[0]	<= 24'b11111110_11111110_11111110; // 白
		RGB_reg	[1]	<= 24'b00000000_11111110_00000000; // 红 
		RGB_reg	[2]	<= 24'b11001101_11111110_00000000; // 橙
		RGB_reg	[3]	<= 24'b11111110_11111110_00000000; // 黄
		RGB_reg	[4]	<= 24'b11111110_00000000_00000000; // 绿
		RGB_reg	[5]	<= 24'b11111110_00000000_11111110; // 青
		RGB_reg	[6]	<= 24'b00000000_00000000_11111110; // 蓝 
		RGB_reg	[7]	<= 24'b00000000_11001100_11001100; // 紫
		RGB_reg	[8]	<= 24'b00000000_00000000_00000000;
		end
		
		10'b0000010000 :  begin
	  	RGB_reg	[0]	<= 24'b00000000_11001100_11001100; // 紫
		RGB_reg	[1]	<= 24'b11111110_11111110_11111110; // 白
		RGB_reg	[2]	<= 24'b00000000_11111110_00000000; // 红
		RGB_reg	[3]	<= 24'b11001101_11111110_00000000; // 橙
		RGB_reg	[4]	<= 24'b11111110_11111110_00000000; // 黄
		RGB_reg	[5]	<= 24'b11111110_00000000_00000000; // 绿
		RGB_reg	[6]	<= 24'b11111110_00000000_11111110; // 青
		RGB_reg	[7]	<= 24'b00000000_00000000_11111110; // 蓝
		RGB_reg	[8]	<= 24'b00000000_00000000_00000000;
		end
		
		10'b0000100000 :  begin
	  	RGB_reg	[0]	<= 24'b00000000_00000000_11111110; // 蓝
		RGB_reg	[1]	<= 24'b00000000_11001100_11001100; // 紫
		RGB_reg	[2]	<= 24'b11111110_11111110_11111110; // 白
		RGB_reg	[3]	<= 24'b00000000_11111110_00000000; // 红
		RGB_reg	[4]	<= 24'b11001101_11111110_00000000; // 橙
		RGB_reg	[5]	<= 24'b11111110_11111110_00000000; // 黄
		RGB_reg	[6]	<= 24'b11111110_00000000_00000000; // 绿
		RGB_reg	[7]	<= 24'b11111110_00000000_11111110; // 青
		RGB_reg	[8]	<= 24'b00000000_00000000_00000000;
		end
		
		10'b0001000000 :  begin
	  	RGB_reg	[0]	<= 24'b11111110_00000000_11111110; // 青
		RGB_reg	[1]	<= 24'b00000000_00000000_11111110; // 蓝
		RGB_reg	[2]	<= 24'b00000000_11001100_11001100; // 紫
		RGB_reg	[3]	<= 24'b11111110_11111110_11111110; // 白
		RGB_reg	[4]	<= 24'b00000000_11111110_00000000; // 红
		RGB_reg	[5]	<= 24'b11001101_11111110_00000000; // 橙
		RGB_reg	[6]	<= 24'b11111110_11111110_00000000; // 黄
		RGB_reg	[7]	<= 24'b11111110_00000000_00000000; // 绿
		RGB_reg	[8]	<= 24'b00000000_00000000_00000000;
		end
		
		10'b0010000000 :  begin
	  	RGB_reg	[0]	<= 24'b11111110_00000000_00000000; // 绿
		RGB_reg	[1]	<= 24'b11111110_00000000_11111110; // 青
		RGB_reg	[2]	<= 24'b00000000_00000000_11111110; // 蓝
		RGB_reg	[3]	<= 24'b00000000_11001100_11001100; // 紫
		RGB_reg	[4]	<= 24'b11111110_11111110_11111110; // 白
		RGB_reg	[5]	<= 24'b00000000_11111110_00000000; // 红
		RGB_reg	[6]	<= 24'b11001101_11111110_00000000; // 橙
		RGB_reg	[7]	<= 24'b11111110_11111110_00000000; // 黄
		RGB_reg	[8]	<= 24'b00000000_00000000_00000000;
		end
		
		10'b0100000000 :  begin
	  	RGB_reg	[0]	<= 24'b11111110_11111110_00000000; // 黄
		RGB_reg	[1]	<= 24'b11111110_00000000_00000000; // 绿
		RGB_reg	[2]	<= 24'b11111110_00000000_11111110; // 青
		RGB_reg	[3]	<= 24'b00000000_00000000_11111110; // 蓝
		RGB_reg	[4]	<= 24'b00000000_11001100_11001100; // 紫
		RGB_reg	[5]	<= 24'b11111110_11111110_11111110; // 白
		RGB_reg	[6]	<= 24'b00000000_11111110_00000000; // 红
		RGB_reg	[7]	<= 24'b11001101_11111110_00000000; // 橙
		RGB_reg	[8]	<= 24'b00000000_00000000_00000000;
		end
		
		10'b1000000000 :  begin
	  	RGB_reg	[0]	<= 24'b11001101_11111110_00000000; // 橙
		RGB_reg	[1]	<= 24'b11111110_11111110_00000000; // 黄
		RGB_reg	[2]	<= 24'b11111110_00000000_00000000; // 绿
		RGB_reg	[3]	<= 24'b11111110_00000000_11111110; // 青
		RGB_reg	[4]	<= 24'b00000000_00000000_11111110; // 蓝
		RGB_reg	[5]	<= 24'b00000000_11001100_11001100; // 紫
		RGB_reg	[6]	<= 24'b11111110_11111110_11111110; // 白
		RGB_reg	[7]	<= 24'b00000000_11111110_00000000; // 红
		RGB_reg	[8]	<= 24'b00000000_00000000_00000000;
		end
		endcase
	end
	else if(uart_data[6]) begin   
//3. 闪烁+红绿蓝白移位循环
	case(mode)    
	   10'b0000000001 :  begin
	   RGB_reg	[0]	<= 24'b00000000_11111110_00000000; // 红
		RGB_reg	[1]	<= 24'b11001101_11111110_00000000; // 橙
		RGB_reg	[2]	<= 24'b11111110_11111110_00000000; // 黄
		RGB_reg	[3]	<= 24'b11111110_00000000_00000000; // 绿
		RGB_reg	[4]	<= 24'b11111110_00000000_11111110; // 青
		RGB_reg	[5]	<= 24'b00000000_00000000_11111110; // 蓝
		RGB_reg	[6]	<= 24'b00000000_11001100_11001100; // 紫
		RGB_reg	[7]	<= 24'b11111110_11111110_11111110; // 白
		RGB_reg	[8]	<= 24'b11111111_11111111_11111111;
		end

      10'b0000000010 :  begin
	  	RGB_reg	[0]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[1]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[2]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[3]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[4]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[5]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[6]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[7]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[8]	<= 24'b00000000_00000000_00000000;
		end

      //红绿蓝白红绿蓝白循环
		10'b0000000100 :  begin
	  	RGB_reg	[0]	<= 24'b00000000_11111110_00000000; 
		RGB_reg	[1]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[2]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[3]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[4]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[5]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[6]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[7]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[8]	<= 24'b00000000_00000000_00000000;
		end
		
		10'b0000001000 :  begin
	  	RGB_reg	[0]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[1]	<= 24'b11111110_00000000_00000000;  
		RGB_reg	[2]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[3]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[4]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[5]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[6]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[7]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[8]	<= 24'b00000000_00000000_00000000;
		end
		
		10'b0000010000 :  begin
	  	RGB_reg	[0]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[1]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[2]	<= 24'b00000000_00000000_11111110;  
		RGB_reg	[3]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[4]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[5]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[6]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[7]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[8]	<= 24'b00000000_00000000_00000000;
		end
		
		10'b0000100000 :  begin
	  	RGB_reg	[0]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[1]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[2]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[3]	<= 24'b11111110_11111110_11111110;  
		RGB_reg	[4]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[5]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[6]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[7]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[8]	<= 24'b00000000_00000000_00000000;
		end
		
		10'b0001000000 :  begin
	  	RGB_reg	[0]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[1]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[2]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[3]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[4]	<= 24'b00000000_11111110_00000000; 
		RGB_reg	[5]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[6]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[7]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[8]	<= 24'b00000000_00000000_00000000;
		end
		
		10'b0010000000 :  begin
	  	RGB_reg	[0]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[1]	<= 24'b00000000_00000000_00000000;  
		RGB_reg	[2]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[3]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[4]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[5]	<= 24'b11111110_00000000_00000000; 
		RGB_reg	[6]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[7]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[8]	<= 24'b00000000_00000000_00000000;
		end
		
		10'b0100000000 :  begin
	  	RGB_reg	[0]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[1]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[2]	<= 24'b00000000_00000000_00000000;  
		RGB_reg	[3]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[4]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[5]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[6]	<= 24'b00000000_00000000_11111110; 
		RGB_reg	[7]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[8]	<= 24'b00000000_00000000_00000000;
		end
		
		10'b1000000000 :  begin
	  	RGB_reg	[0]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[1]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[2]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[3]	<= 24'b00000000_00000000_00000000;  
		RGB_reg	[4]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[5]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[6]	<= 24'b00000000_00000000_00000000; 
		RGB_reg	[7]	<= 24'b11111110_11111110_11111110; 
		RGB_reg	[8]	<= 24'b00000000_00000000_00000000;
		end
		endcase
	end
	else if(uart_data[7]) begin   
//4. 全亮
	case(mode)    
	   10'b0000000001 :  begin
	   RGB_reg	[0]	<= 24'b00011111_00011111_00011111; // 红
		RGB_reg	[1]	<= 24'b00011111_00011111_00011111; // 橙
		RGB_reg	[2]	<= 24'b00011111_00011111_00011111; // 黄
		RGB_reg	[3]	<= 24'b00011111_00011111_00011111; // 绿
		RGB_reg	[4]	<= 24'b00011111_00011111_00011111; // 青
		RGB_reg	[5]	<= 24'b00011111_00011111_00011111; // 蓝
		RGB_reg	[6]	<= 24'b00011111_00011111_00011111; // 紫
		RGB_reg	[7]	<= 24'b00011111_00011111_00011111; // 白
		RGB_reg	[8]	<= 24'b00011111_00011111_00011111;
		end

      10'b0000000010 :  begin
	  	RGB_reg	[0]	<= 24'b00011111_00011111_00011111; 
		RGB_reg	[1]	<= 24'b00011111_00011111_00011111; 
		RGB_reg	[2]	<= 24'b00011111_00011111_00011111; 
		RGB_reg	[3]	<= 24'b00011111_00011111_00011111; 
		RGB_reg	[4]	<= 24'b00011111_00011111_00011111; 
		RGB_reg	[5]	<= 24'b00011111_00011111_00011111; 
		RGB_reg	[6]	<= 24'b00011111_00011111_00011111; 
		RGB_reg	[7]	<= 24'b00011111_00011111_00011111; 
		RGB_reg	[8]	<= 24'b00011111_00011111_00011111;
		end

      //红绿蓝白红绿蓝白循环
		10'b0000000100 :  begin
	  	RGB_reg	[0]	<= 24'b00011111_00011111_00011111; 
		RGB_reg	[1]	<= 24'b00011111_00011111_00011111; 
		RGB_reg	[2]	<= 24'b00011111_00011111_00011111; 
		RGB_reg	[3]	<= 24'b00011111_00011111_00011111; 
		RGB_reg	[4]	<= 24'b00011111_00011111_00011111; 
		RGB_reg	[5]	<= 24'b00011111_00011111_00011111; 
		RGB_reg	[6]	<= 24'b00011111_00011111_00011111; 
		RGB_reg	[7]	<= 24'b00011111_00011111_00011111; 
		RGB_reg	[8]	<= 24'b00011111_00011111_00011111;
		end
		
		10'b0000001000 :  begin
	  	RGB_reg	[0]	<= 24'b00011111_00011111_00011111; 
		RGB_reg	[1]	<= 24'b00011111_00011111_00011111;  
		RGB_reg	[2]	<= 24'b00011111_00011111_00011111; 
		RGB_reg	[3]	<= 24'b00011111_00011111_00011111; 
		RGB_reg	[4]	<= 24'b00011111_00011111_00011111; 
		RGB_reg	[5]	<= 24'b00011111_00011111_00011111; 
		RGB_reg	[6]	<= 24'b00011111_00011111_00011111; 
		RGB_reg	[7]	<= 24'b00011111_00011111_00011111; 
		RGB_reg	[8]	<= 24'b00011111_00011111_00011111;
		end
		
		10'b0000010000 :  begin
	  	RGB_reg	[0]	<= 24'b00011111_00011111_00011111; 
		RGB_reg	[1]	<= 24'b00011111_00011111_00011111; 
		RGB_reg	[2]	<= 24'b00011111_00011111_00011111;  
		RGB_reg	[3]	<= 24'b00011111_00011111_00011111; 
		RGB_reg	[4]	<= 24'b00011111_00011111_00011111; 
		RGB_reg	[5]	<= 24'b00011111_00011111_00011111; 
		RGB_reg	[6]	<= 24'b00011111_00011111_00011111; 
		RGB_reg	[7]	<= 24'b00011111_00011111_00011111; 
		RGB_reg	[8]	<= 24'b00011111_00011111_00011111;
		end
		
		10'b0000100000 :  begin
	  	RGB_reg	[0]	<= 24'b00011111_00011111_00011111; 
		RGB_reg	[1]	<= 24'b00011111_00011111_00011111; 
		RGB_reg	[2]	<= 24'b00011111_00011111_00011111; 
		RGB_reg	[3]	<= 24'b00011111_00011111_00011111;  
		RGB_reg	[4]	<= 24'b00011111_00011111_00011111; 
		RGB_reg	[5]	<= 24'b00011111_00011111_00011111; 
		RGB_reg	[6]	<= 24'b00011111_00011111_00011111; 
		RGB_reg	[7]	<= 24'b00011111_00011111_00011111; 
		RGB_reg	[8]	<= 24'b00011111_00011111_00011111;
		end
		
		10'b0001000000 :  begin
	  	RGB_reg	[0]	<= 24'b00011111_00011111_00011111; 
		RGB_reg	[1]	<= 24'b00011111_00011111_00011111; 
		RGB_reg	[2]	<= 24'b00011111_00011111_00011111; 
		RGB_reg	[3]	<= 24'b00011111_00011111_00011111; 
		RGB_reg	[4]	<= 24'b00011111_00011111_00011111; 
		RGB_reg	[5]	<= 24'b00011111_00011111_00011111; 
		RGB_reg	[6]	<= 24'b00011111_00011111_00011111; 
		RGB_reg	[7]	<= 24'b00011111_00011111_00011111; 
		RGB_reg	[8]	<= 24'b00011111_00011111_00011111;
		end
		
		10'b0010000000 :  begin
	  	RGB_reg	[0]	<= 24'b00011111_00011111_00011111; 
		RGB_reg	[1]	<= 24'b00011111_00011111_00011111;  
		RGB_reg	[2]	<= 24'b00011111_00011111_00011111; 
		RGB_reg	[3]	<= 24'b00011111_00011111_00011111; 
		RGB_reg	[4]	<= 24'b00011111_00011111_00011111; 
		RGB_reg	[5]	<= 24'b00011111_00011111_00011111; 
		RGB_reg	[6]	<= 24'b00011111_00011111_00011111; 
		RGB_reg	[7]	<= 24'b00011111_00011111_00011111; 
		RGB_reg	[8]	<= 24'b00011111_00011111_00011111;
		end
		
		10'b0100000000 :  begin
	  	RGB_reg	[0]	<= 24'b00011111_00011111_00011111; 
		RGB_reg	[1]	<= 24'b00011111_00011111_00011111; 
		RGB_reg	[2]	<= 24'b00011111_00011111_00011111;  
		RGB_reg	[3]	<= 24'b00011111_00011111_00011111; 
		RGB_reg	[4]	<= 24'b00011111_00011111_00011111; 
		RGB_reg	[5]	<= 24'b00011111_00011111_00011111; 
		RGB_reg	[6]	<= 24'b00011111_00011111_00011111; 
		RGB_reg	[7]	<= 24'b00011111_00011111_00011111; 
		RGB_reg	[8]	<= 24'b00011111_00011111_00011111;
		end
		
		10'b1000000000 :  begin
	  	RGB_reg	[0]	<= 24'b00011111_00011111_00011111; 
		RGB_reg	[1]	<= 24'b00011111_00011111_00011111; 
		RGB_reg	[2]	<= 24'b00011111_00011111_00011111; 
		RGB_reg	[3]	<= 24'b00011111_00011111_00011111;  
		RGB_reg	[4]	<= 24'b00011111_00011111_00011111; 
		RGB_reg	[5]	<= 24'b00011111_00011111_00011111; 
		RGB_reg	[6]	<= 24'b00011111_00011111_00011111; 
		RGB_reg	[7]	<= 24'b00011111_00011111_00011111; 
		RGB_reg	[8]	<= 24'b00011111_00011111_00011111;
		end
		endcase
	end
end

//===============================================//
//===================================================//

always @(posedge clk_RGB_Control or negedge rst_n) begin
	if(!rst_n)	begin
		k <= 0;
		RGB <= 0;
	end
	else if(tx_en_r)	begin    //tx_en_r发送数据控制使能
		case (k)
			5'd0,5'd1,5'd2,5'd3,5'd4,5'd5,5'd6,5'd7:
				if(tx_done_r0)	begin
					RGB <= RGB_reg[k];
					k <= k + 1;
				end
			5'd8:
				if(tx_done)	begin
					RGB <= RGB_reg[0];
					k <= 0;
				end
		  	default: k <= 0;
		endcase
	end
	else ;
end
//--------------------------------//

//-------------计数器-------------//
always @(posedge clk_RGB_Control) begin
	if((!rst_n) || (tx_en_r))	begin  //tx_en_r发送数据控制使能
		cnt <= 0;
	end
	else if(cnt == 32'd14999)	begin	//RESET时间(300us*50M=15000)
		cnt <= cnt;
	end
	else	begin
		cnt <= cnt + 1;
	end
end
//--------------------------------//

//--------------------------------//
always @(posedge clk_RGB_Control or negedge rst_n) begin   //tx_en_r 发送数据控制使能
	if(!rst_n)	begin
		tx_en_r <= 0;
	end
	else if((k == 5'd8) && (tx_done))	begin
		tx_en_r <= 0;			//一组数据发送结束，RESTE
	end
	else if((cnt == 32'd14999) && tx_done)	begin
		tx_en_r <= 1;			//重新开始发送
	end
	else	begin
		tx_en_r <= tx_en_r;
	end
end

assign	tx_en = tx_en_r;
//--------------------------------//
endmodule
