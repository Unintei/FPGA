/*****************************************************

*****************************************************/
module  SUM_Led
#(
//****************************************************//

//定义晶振频率50M
    parameter Red = 3'b011  ,

    parameter Yellow = 3'b101,

    parameter Green = 3'b110 
	
//****************************************************//
)
(
    input   wire            sys_clk     ,   //输入工作时钟,频率50MHz
    input   wire            sys_rst_n   ,   //输入复位信号,低电平有效

	output  wire    [3:0]    sum_cnt		,
    output  wire    [6:0]    sum_out         ,
	output  wire    [2:0]    Led		,
	
	output  wire    [2:0]    Led2		
);

wire     [ 5:0]  cnt1         ;    //0.1ms
wire     [ 5:0]  x1         ;    //0.1ms

wire     [ 5:0]  cnt2         ;    //0.1ms
wire     [ 5:0]  x2         ;    //0.1ms
//********************************************************************//
//***************************** Main Code ****************************//
//********************************************************************//
//***************************** Main Code ****************************//
//********************************************************************//
//***************************** Main Code ****************************//
//********************************************************************//

led  led1(
		.sys_clk  	(sys_clk)  ,   //输入工作时钟,频率50MHz
		.sys_rst_n	(sys_rst_n)  ,   //输入复位信号,低电平有效
		.sel		(Yellow)    ,

		.x			(x1),

		.cnt2		(cnt1),
		.led_sel  	(Led)
);


led  led2(
		.sys_clk  	(sys_clk)  ,   //输入工作时钟,频率50MHz
		.sys_rst_n	(sys_rst_n)  ,   //输入复位信号,低电平有效
		.sel		(Red)    ,

		.x			(x2),

		.cnt2		(cnt2),
		.led_sel  	(Led2)
);

sum  sum(
		.sys_clk	(sys_clk)  ,   //输入工作时钟,频率50MHz
		.sys_rst_n	(sys_rst_n)  ,   //输入复位信号,低电平有效
		
		.cnt1		(cnt1),
		.x1			(x1),

		.cnt2		(cnt2),
		.x2			(x2),
		
		.seg_sel	(sum_cnt),
		.seg_ment	(sum_out)
);

endmodule
