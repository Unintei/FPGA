/*****************************************************
	动态数码管 
	2023/11/21    1s切换一位
*****************************************************/
module  SUM_Led
#(
//****************************************************//

//定义晶振频率50M
    parameter CNT_MAX = 26'd50_000_000 
	 
//****************************************************//
)
(
    input   wire            sys_clk     ,   //输入工作时钟,频率50MHz
    input   wire            sys_rst_n   ,   //输入复位信号,低电平有效

	 output  wire    [7:0]    Led_cnt		,
    output  wire    [6:0]    led          //输出行同步信号

);


wire end_cnt0 ;

//********************************************************************//
//***************************** Main Code ****************************//
//********************************************************************//

  jsq jsq1
(
   .sys_clk  (sys_clk)   ,   //输入工作时钟,频率50MHz
   .sys_rst_n(sys_rst_n)   ,   //输入复位信号,低电平有效
	
   .end_cnt0 (end_cnt0)         //输出行同步信号

);

//********************************************************************//
//***************************** Main Code ****************************//
//********************************************************************//

  cen cen1
(
    .sys_clk    (sys_clk) ,   //输入工作时钟,频率50MHz
    .sys_rst_n  (sys_rst_n) ,   //输入复位信号,低电平有效
    .end_cnt0   (end_cnt0) ,
					
	.Led_cnt	(Led_cnt)	

);

//********************************************************************//
//***************************** Main Code ****************************//
//********************************************************************//
ymq ymq1
(
	.sys_clk    (sys_clk),
	.sys_rst_n  (sys_rst_n),
	.Led_cnt	(Led_cnt),
	.end_cnt0(end_cnt0),
   .led		(led)       

);

endmodule
