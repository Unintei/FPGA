/*****************************************************
	动态数码管 
	2023/11/21    1s切换一位
*****************************************************/
module  cen
#(
//****************************************************//

//定义晶振频率50M
    parameter CNT_MAX = 26'd50_000_000 
	 
//****************************************************//
)
(
    input   wire            sys_clk     ,   //输入工作时钟,频率50MHz
    input   wire            sys_rst_n   ,   //输入复位信号,低电平有效
    input   wire            end_cnt0    ,

	output  reg    [7:0]    Led_cnt		

);






//********************************************************************//
//***************************** Main Code ****************************//
//********************************************************************//

//Led_cnt:数码管片选信号
always @(posedge sys_clk or negedge sys_rst_n)begin
    if(!sys_rst_n)begin  
        Led_cnt <= 8'b1111_1110;
    end
    else if(end_cnt0)	//1s到了
	
            Led_cnt <={Led_cnt[6:0],Led_cnt[7]};   
		 else
            Led_cnt <= Led_cnt;
end


endmodule
